module bcd_gate(a, y);

    input [3:0] a;
    output reg [6:0] y;

    always @(a) begin
        case (a)
            4'b0000: y = 7'b1111110; //0
            4'b0001: y = 7'b0110000; //1
            4'b0010: y = 7'b1101101; //2
            4'b0011: y = 7'b1111001; //3
            4'b0100: y = 7'b0110011; //4
            4'b0101: y = 7'b1011011; //5
            4'b0110: y = 7'b1011111; //6
            4'b0111: y = 7'b1110000; //7
            4'b1000: y = 7'b1111111; //8
            4'b1001: y = 7'b1111011; //9
            4'b1010: y = 7'b1110111; //A
            4'b1011: y = 7'b0011111; //B
            4'b1100: y = 7'b1001110; //C
            4'b1101: y = 7'b0111101; //D
            4'b1110: y = 7'b1001111; //E
            4'b1111: y = 7'b1000111; //F
            default: y = 7'b0000000;
        endcase
    end

endmodule